.PARAM
+ LM1 = 5.0945e-07
+ LM2 = 7.2333e-07
+ LM3 = 1.0093e-06
+ WM1 = 8.8127e-05
+ WM2 = 7.5044e-05
+ WM3 = 9.6361e-06
+ Ib = 0.00012374
