.PARAM
+ LM1 = 4.4703e-07
+ LM2 = 5.6229e-07
+ LM3 = 1.0502e-06
+ WM1 = 8.9235e-05
+ WM2 = 6.7093e-05
+ WM3 = 1.2311e-05
+ Ib = 0.00028325
