.PARAM
+ LM1 = 4.7572e-07
+ LM2 = 4.2032e-07
+ LM3 = 9.2271e-07
+ WM1 = 8.7781e-05
+ WM2 = 7.3793e-05
+ WM3 = 1.1604e-05
+ Ib = 0.00013385
