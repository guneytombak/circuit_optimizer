.PARAM
+ LM1 = 2.2929e-07
+ LM2 = 4.6526e-07
+ LM3 = 4.2452e-07
+ WM1 = 7.9593e-05
+ WM2 = 7.2058e-05
+ WM3 = 2.4235e-05
+ Ib = 0.00028014
