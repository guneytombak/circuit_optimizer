.PARAM
+ WM1 = 8.8365e-05
+ WM2 = 5.3811e-05
+ WM3 = 6.5978e-05
+ WM4 = 0.0001444
+ WM5 = 0.00012508
+ WM6 = 0.00011073
+ WM7 = 4.4437e-05
+ WM8 = 6.8879e-05
+ WM9 = 0.00013067
+ WM10 = 0.00010566
+ WM11 = 3.1785e-05
+ Lcm = 1.2185e-06
+ Rb = 20013.718
+ Cff = 5.3255e-12
